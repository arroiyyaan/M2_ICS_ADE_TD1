library ieee;
use ieee.std_logic_1164.all;
entity test_exemple is
	-- Empty entity
end entity test_exemple;
