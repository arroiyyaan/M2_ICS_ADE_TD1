library ieee;
use ieee.std_logic_1164.all;
entity example is
	port (
		a : in std_logic;
		b : in std_logic;
		c : in std_logic;bluet	
		s1 : out std_logic;
		s2 : out std_logic
	);
end entity example;
